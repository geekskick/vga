library ieee;
use ieee.std_logic_1164.all;

entity top_vga_tb is
end top_vga_tb;

architecture Behavioral of top_vga_tb is   
begin
end Behavioral;